-- EJEMPLO CODIGO MULIPLEXOR 2 A 1 VHDL
-- MUX.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX IS 
PORT (I: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
A,B: IN STD_LOGIC;
Q: OUT STD_LOGIC);
END MUX;

ARCHITECTURE BETTER OF MUX IS 
BEGIN 
PROCESS (I, A, B)
VARIABLE MUXVAL : INTEGER;
BEGIN 
MUXVAL := 0;                                -- ASIGNACION IMPLICITA
IF (A = '1') THEN 
MUXVAL := MUXVAL + 1;
END IF;

IF (b = '1') THEN 
MUXVAL := MUXVAL + 1;
END IF; 

CASE MUXVAL IS                              -- CASE VARIABLE IS ... 
WHEN 0 =>
Q <= IO(0) AFTER 10 NS;
WHEN 1 =>
Q <= IO(1) AFTER 10 NS;
WHEN 2 =>
Q <= IO(2) AFTER 10 NS; 
WHEN 3 =>
Q <= IO(3) AFTER 10 NS;
WHEN OTHERS => 
NULL;
END CASE; 
END PROCESS;
END BETTER;