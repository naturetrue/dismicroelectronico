LIBRARY IEEE;
USE IEEE.STD_LOGIC1164.ALL;
PACKAGE SIGDEC1 IS 
TYPE BUS_TYPE IS ARRAY (0 TO 7) OF STD_LOGIC;

SIGNAL VCC : STD_LOGIC := '1';
SIGNAL GND : STD_LOGIC := '0';

FUNCTION MAGIC_FUNCTION(A : IN BUS_TYPE) RETURN BUS_TYPE;
END SIGNAL;

USE WORK.SIGDEC.ALL;
LIBRARY IEEE;
 
---------------------------------------------------------

UNSIGNED 
INTEGER 
SIGNED 
STD_LOGIC_VECTOR
STD_LOGIC 
BIT 
BIT_VECTOR 
