-- EJEMPLO ASIGNACIONES SECUENCIALES
-- NAND2.VHD

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY NAND2 IS 
PORT(A,B : IN STD_LOGIC;
C : OUT STD_LOGIC);
END NAND2;

ARCHITECTURE NAND2 OF NAND2 IS  -- FORMULACION DE UN ARCHITECTURE --> ARCHITECTURE NOMBRE_ARCH OF NOMBRE_ENT IS
BEGIN 
PROCESS (a, B)                  -- SENALES A LAS QUE RESPONDE 
VARIABLE TEMP : STD_LOGIC;      -- VARIABLES EN VHDL (SE LES PUEDE ASIGNAR VALORES DE FORMA DINAMICA), DE FORMA ESTATICA USAR CONSTANT
BEGIN 
TEMP := NOT (A AND B);
IF (TEMP = '1') THEN 
C <= TEMP AFTER 6 NS; 
ELSIF (TEMP = '0') THEN 
C <= TEMP AFTER 5 NS;
ELSE 
C <= TEMP AFTER 6 NS; 
END IF ;
END PROCESS;
END NAND2;