LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY TEST IS 
GENERIC (RISE, FALL : TIME;
LOAD : INTEGER);
PORT (INA, INB,INC,IND: IN STD_LOGIC;
OUT1,OUT2: OUT STD_LOGIC);
END TEST;

ARCHITECTURE TEST_ARCH OF TEST IS 
COMPONENT AND2
GENERIC(RISE,FALL: TIME := 10 NS;
LOAD : INTEGER := 0);
PORT(A,B:IN STD_LOGIC;
C:OUT STD_LOGIC);
END COMPONENT;
BEGIN 
U1: AND2 GENERIC MAP (10 NS,12 NS, 3)
PORT MAP (INA, INB, INC);
U2: AND2 PORT MAP (INC, IND, OUT2);
END TEST_ARCH;
